.model MYSW SW(Ron=1 Roff=1Meg Vt=.5 Vh=-.4)
